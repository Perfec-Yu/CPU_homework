module WB();
	// deleted
endmodule
